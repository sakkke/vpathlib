module vpathlib
